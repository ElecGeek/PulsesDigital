library ieee;
use ieee.std_logic_1164.all;

entity Amplitudes_multiplier_test is

end entity Amplitudes_multiplier_test;

architecture arch of Amplitudes_multiplier_test is

begin

end architecture arch;
